// Jason Bowman
// jbowman@hmc.edu
// CREATED: 10-28-24
// This module acts as the add round key part of AES, using XOR with the appropriate input depending on the round and throwing a flag once each round has been completed

